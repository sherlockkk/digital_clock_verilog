module print2(fs,a,b,c,d,e,f,led_dig,display);
input fs;
input [3:0]a,b,c,d,e,f;

output [7:0]led_dig,display;
reg	   [7:0]led_dig,display;

reg    [3:0]o;
always @(posedge fs)
begin
    case(o)
		4'b0000:begin
					led_dig<=8'b11101111;
			          case(a)//1/100���λѡ����ʾ
			              4'b0000:begin display<=8'b0111111;end
			              4'b0001:begin display<=8'b0000110;end
			              4'b0010:begin display<=8'b1011011;end
			              4'b0011:begin display<=8'b1001111;end
			              4'b0100:begin display<=8'b1100110;end
			              4'b0101:begin display<=8'b1101101;end
			              4'b0110:begin display<=8'b1111101;end
			              4'b0111:begin display<=8'b0000111;end
			              4'b1000:begin display<=8'b1111111;end
			              4'b1001:begin display<=8'b1101111;end
			              default:;
				 	 endcase
       			end
       4'b0001:begin
				led_dig<=8'b11110111;
					   case(b)//1/100���λѡ����ʾ
			              4'b0000:begin display<=8'b0111111;end
			              4'b0001:begin display<=8'b0000110;end
			              4'b0010:begin display<=8'b1011011;end
			              4'b0011:begin display<=8'b1001111;end
			              4'b0100:begin display<=8'b1100110;end
			              4'b0101:begin display<=8'b1101101;end
				      4'b0110:begin display<=8'b1111101;end
			              4'b0111:begin display<=8'b0000111;end
			              4'b1000:begin display<=8'b1111111;end
			              4'b1001:begin display<=8'b1101111;end	
			              default:;
		         	 endcase
       			end
		4'b0010: begin led_dig<=8'b11111101;display<=8'b1000000;end
		4'b0011:begin
				led_dig<=8'b11111110;
				   case(c)//���λѡ����ʾ
		              4'b0000:begin display<=8'b0111111;end
		              4'b0001:begin display<=8'b0000110;end
		              4'b0010:begin display<=8'b1011011;end
		              4'b0011:begin display<=8'b1001111;end
		              4'b0100:begin display<=8'b1100110;end
		              4'b0101:begin display<=8'b1101101;end
		              4'b0110:begin display<=8'b1111101;end
		              4'b0111:begin display<=8'b0000111;end
		              4'b1000:begin display<=8'b1111111;end
		              4'b1001:begin display<=8'b1101111;end
						default:;
		          endcase
          		end
      4'b0100:begin
			led_dig<=8'b11111011;
			case(d)//���λѡ����ʾ
	              4'b0000:begin display<=8'b0111111;end
	              4'b0001:begin display<=8'b0000110;end
	              4'b0010:begin display<=8'b1011011;end
	              4'b0011:begin display<=8'b1001111;end
	              4'b0100:begin display<=8'b1100110;end
	              4'b0101:begin display<=8'b1101101;end
	              default:;
	        endcase
       	 end		
		4'b0101: begin led_dig<=8'b01111111;display<=8'b1000000;end
		4'b0110:begin
			   led_dig<=8'b10111111;
				case(e)//�ֵ�λѡ����ʾ
		              4'b0000:begin display<=8'b0111111;end
		              4'b0001:begin display<=8'b0000110;end
		              4'b0010:begin display<=8'b1011011;end
		              4'b0011:begin display<=8'b1001111;end
		              4'b0100:begin display<=8'b1100110;end
		              4'b0101:begin display<=8'b1101101;end
		              4'b0110:begin display<=8'b1111101;end
		              4'b0111:begin display<=8'b0000111;end
		              4'b1000:begin display<=8'b1111111;end
		              4'b1001:begin display<=8'b1101111;end
						default:;
			  	endcase             
       			end
		4'b0111:begin
				led_dig<=8'b11011111;
				   case(f)//�ָ�λѡ����ʾ
		              4'b0000:begin display<=8'b0111111;end
		              4'b0001:begin display<=8'b0000110;end
		              4'b0010:begin display<=8'b1011011;end
		              default:;
		          endcase
	      		end
		default:;
		endcase
	o<=o+4'b0001;
	if(o===4'b0111)o<=4'b0000;	
end//������ʱ����
endmodule